`ifndef DEFS_SVH
`define DEFS_SVH
`define CACHE_SIZE 4096
`define CACHE_BLOCKS 256
`define CACHE_LINE_SIZE 128
`define CACHE_TAG_SIZE 20
`define OPCODE_L 2
`define OPCODE_S 3
`endif // DEFS_SVH


