`ifndef array_mul
`define array_mul

parameter width = 16;
parameter result_width = 32;

`endif