`ifndef restor_div
`define restor_div

parameter  width = 32;
parameter  counter_width = 5;

`endif 