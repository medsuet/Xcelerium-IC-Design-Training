module tb_sequential_adder;

    // Testbench signals
    logic clk;
    logic reset;
    logic [3:0] number;
    logic output_lsb;

    // Instantiate the design under test (DUT)
    sequential_adder dut (
        .clk(clk),
        .reset(reset),
        .number(number),
        .output_lsb(output_lsb)
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 10ns period clock
    end

    // Task to apply reset
    task apply_reset();
        begin
            @(posedge clk);
            reset = 1;
            @(posedge clk);
            reset = 0;
        end
    endtask

    // Task to apply a test case
    task apply_test_case(input logic [3:0] test_number);
        begin
            number = test_number;
            repeat(4) @(posedge clk);  // Wait enough time for the FSM to process the number
        end
    endtask

    // Test sequence
    initial begin
        // Initialize signals
        clk = 0;
        reset = 0;
        number = 4'b0000;

        // Apply reset
        apply_reset();

        // Apply test cases using a for loop
        for (int i = 0; i < 16; i++) begin
            apply_test_case(i[3:0]);
        end

        // End of simulation
        $finish;
    end

    // Monitor the output
    initial begin
        $monitor("Time: %0t, Reset: %b, Number: %b, Output LSB: %b", $time, reset, number, output_lsb);
    end

    // Generate VCD file for waveform analysis
    initial begin
        $dumpfile("sequential_adder.vcd");
        $dumpvars(0, tb_sequential_adder);
    end

endmodule
