module tb_restoring_division;
endmodule