/*
    Name: SequentialSignedMultiplier.sv
    Author: Muhammad Tayyab
    Date: 30-7-2024
    Description: Testbench for SequentialSignedMultiplier.sv
*/

//`define DIRECTEDTEST

module SequentialSignedMultiplier_tb();
    parameter NUMTESTS = 1e1;
    parameter NUMBITS = 16;
int i;
    logic clk, reset, start;
    logic [(NUMBITS-1):0] numA, numB;
    logic ready;
    logic [((2*NUMBITS)-1):0] test_result, ref_result;

    SequentialSignedMultiplier #(NUMBITS) ssm
    (
        clk, reset, start,
        numA, numB,
        ready,
        test_result
    );

    initial begin
        clk = 1;
        forever #5 clk = ~clk;
    end

    // Directed tests
    `ifdef DIRECTEDTEST
        initial begin
            directed_test(54793,22115);
            directed_test(-1,2);
        end
    `endif

    // Random tests
    `ifndef DIRECTEDTEST
        initial driver();
        initial monitor();
    `endif

    task directed_test(shortint a, shortint b);
        reset_sequence();

        numA = a;
        numB = b;
        start_signal();
        
        ref_result = $signed(int'($signed(numA)) * int'($signed(numB)));   

        @(posedge ready);
        if (ref_result !== test_result) begin
            $display("\n\nDirected test failed.\n");
            $display("numA = %d \nnumB = %d", numA, numB);
            $display("Test_result = h'%x", test_result);
            $display("Correct_result = h'%x\n\n", ref_result);
        end
        else begin
            $display("\n\nDirected test on %d * %d passed.\n\n", numA, numB);
        end
        @(posedge clk);
        $stop();

    endtask

    task driver();
        reset_sequence();

        for (i=0; i<NUMTESTS; i++)
        begin
            numA = $random();
            numB = $random();
            start_signal();
            @(posedge ready);
            @(negedge ready);
        end

        $display("\n\nAll %d tests passed.\n\n", NUMTESTS);
        $stop();
    endtask

    task monitor();
        @(negedge reset);
        @(posedge reset);
        forever begin
            @(posedge clk);

            @(posedge ready);
            ref_result = $signed(int'($signed(numA)) * int'($signed(numB)));
            if (ref_result !== test_result) begin
                $display("\n\nTest failed.\n");
                $display("%d, %d", numA, numB);
                $display("\n\nTest_result = h'%x", test_result);
                $display("Correct_result = h'%x\n\n", ref_result);
                $stop();
            end
        end
    endtask

    task reset_sequence();
        reset = 1;
        #3 reset = 0;
        #14 reset = 1;
    endtask

    task start_signal();
        start = 1;
        @(posedge clk);
        start = 0;
    endtask 

endmodule
