`define VERILATOR