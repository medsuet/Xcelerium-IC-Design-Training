`ifndef sig_mul
`define sig_mul

parameter  width  = 16;
parameter result_width = 32;

`endif 