`define VERILATOR
